$display("Hello, World!");
