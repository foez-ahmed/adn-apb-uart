`define DEFAULT_ADDR_WIDTH 5
`define DEFAULT_DATA_WIDTH 32
