module hello_world;

  initial begin
    `include "dummy.svh"
    $finish;
  end

endmodule
